module counternonrecycling_tb;
	
endmodule